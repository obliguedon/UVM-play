module dut (
    dut_if _if
);
    hello_world my_dut();
endmodule
